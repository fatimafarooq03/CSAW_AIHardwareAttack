`timescale 1ns / 1ps  // Corrected syntax

module riscv_core_tb;

// Clock and Reset Signals
reg clk_i;
reg rst_i;

// Memory Signals
reg [31:0] mem_d_data_rd_i;
reg mem_d_accept_i;
reg mem_d_ack_i;
reg mem_d_error_i;
reg [10:0] mem_d_resp_tag_i;
reg mem_i_accept_i;
reg mem_i_valid_i;
reg mem_i_error_i;
reg [31:0] mem_i_inst_i;
reg intr_i;
reg [31:0] reset_vector_i;
reg [31:0] cpu_id_i;

wire [31:0] mem_d_addr_o;
wire [31:0] mem_d_data_wr_o;
wire mem_d_rd_o;
wire [3:0] mem_d_wr_o;
wire mem_d_cacheable_o;
wire [10:0] mem_d_req_tag_o;
wire mem_d_invalidate_o;
wire mem_d_writeback_o;
wire mem_d_flush_o;
wire mem_i_rd_o;
wire mem_i_flush_o;
wire mem_i_invalidate_o;
wire [31:0] mem_i_pc_o;

// Parameters
parameter MEM_CACHE_ADDR_MIN = 32'h80000000;
parameter MEM_CACHE_ADDR_MAX = 32'h8fffffff;

// Instantiate the RISC-V core
riscv_core uut (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .mem_d_data_rd_i(mem_d_data_rd_i),
    .mem_d_accept_i(mem_d_accept_i),
    .mem_d_ack_i(mem_d_ack_i),
    .mem_d_error_i(mem_d_error_i),
    .mem_d_resp_tag_i(mem_d_resp_tag_i),
    .mem_i_accept_i(mem_i_accept_i),
    .mem_i_valid_i(mem_i_valid_i),
    .mem_i_error_i(mem_i_error_i),
    .mem_i_inst_i(mem_i_inst_i),
    .intr_i(intr_i),
    .reset_vector_i(reset_vector_i),
    .cpu_id_i(cpu_id_i),

    .mem_d_addr_o(mem_d_addr_o),
    .mem_d_data_wr_o(mem_d_data_wr_o),
    .mem_d_rd_o(mem_d_rd_o),
    .mem_d_wr_o(mem_d_wr_o),
    .mem_d_cacheable_o(mem_d_cacheable_o),
    .mem_d_req_tag_o(mem_d_req_tag_o),
    .mem_d_invalidate_o(mem_d_invalidate_o),
    .mem_d_writeback_o(mem_d_writeback_o),
    .mem_d_flush_o(mem_d_flush_o),

    .mem_i_rd_o(mem_i_rd_o),
    .mem_i_flush_o(mem_i_flush_o),
    .mem_i_invalidate_o(mem_i_invalidate_o),
    .mem_i_pc_o(mem_i_pc_o)
);

// Clock Generation
always #5 clk_i = ~clk_i;

// Testbench Logic
initial begin
    // Initialize signals
    clk_i = 0;
    rst_i = 1;
    mem_d_data_rd_i = 0;
    mem_d_accept_i = 1;
    mem_d_ack_i = 1;
    mem_d_error_i = 0;
    mem_d_resp_tag_i = 0;
    mem_i_accept_i = 1;
    mem_i_valid_i = 0;
    mem_i_error_i = 0;
    mem_i_inst_i = 32'd0;   // addi/ld
    intr_i = 0;
    reset_vector_i = 32'h80000000;
    cpu_id_i = 0;

    // Apply reset
    repeat (10) begin
      @(posedge clk_i);
    end
    rst_i = 0;

    // Further operations...
    repeat (3) begin
      @(posedge clk_i);
    end
    
    mem_i_inst_i    = 32'b10000000000000000000_01011_0110111;     //LUI  x11, 0x80000
    mem_i_valid_i   = 1'b1;

    @(posedge clk_i);
    mem_i_inst_i    = 32'b10000000000000000000_01011_0110111;     //LUI  x11, 0x80000
    mem_i_valid_i   = 1'b1;

    @(posedge clk_i);
    mem_i_inst_i    = 32'b10010000000000000000_01100_0110111;     //LUI  x12, 0x90000
    mem_i_valid_i   = 1'b1;

    @(posedge clk_i);
    mem_i_inst_i    = 32'b11011110101011011011_01101_0110111;     //LUI  x13, 0xDEADB
    mem_i_valid_i   = 1'b1;

    @(posedge clk_i);
    mem_i_inst_i    = 32'b111011101111_01101_000_01101_0010011;   //ADDI x13, x0,  0xEEF
    mem_i_valid_i   = 1'b1;

    @(posedge clk_i);
    mem_i_valid_i = 1'b0;

    @(posedge clk_i);
    mem_i_inst_i = 32'b0000000_01101_01011_010_00000_0100011;  //SW   x13, x11, 0x0
    mem_i_valid_i = 1'b1;
    $display("[Expectation]At Address=0x80000000, Value=0xdeadaeef is to be written");


    @(posedge clk_i);
    mem_i_inst_i  = 32'b000000000000_00000_000_01110_0010011;   //ADDI x14, x0,  0x0  NOP
    mem_i_valid_i = 1'b1;

    @(posedge clk_i);
    mem_i_inst_i = 32'b0000000_01101_01100_010_00000_0100011;  //SW   x13, x12, 0x0
    mem_i_valid_i = 1'b1;
    $display("[Expectation]At Address=0x90000000, Value=0xdeadaeef is to be written");

    @(posedge clk_i);
    mem_i_inst_i  = 32'b000000000000_00000_000_01110_0010011;   //ADDI x14, x0,  0x0  NOP
    mem_i_valid_i = 1'b1;
end 
    
// Counter for clock cycles
integer cycle_count = 0;

// Add monitor for memory operations and stop the simulation after 50 clock cycles
always @(posedge clk_i) begin
    // Increment the clock cycle counter
    cycle_count = cycle_count + 1;

    // Detect store (SW) operations
    if (|mem_d_wr_o) begin
        $display("[ACTION] At Time=%0t, Address=0x%08x, Value=0x%08x is written", 
                 $time, mem_d_addr_o, mem_d_data_wr_o);
    end

    // Stop the simulation after 50 clock cycles
    if (cycle_count == 50) begin
        //$display("[INFO] Simulation ended after %0d clock cycles.", cycle_count);
        $finish; // End the simulation
    end
end

endmodule
 